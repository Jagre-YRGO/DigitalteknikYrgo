library IEEE;
use IEEE.std_logic_1164.all;

entity spi_slave is
   port
   (
      sclk : in std_logic;
      mosi : in std_logic
   );
end entity;

architecture rtl of spi_slave is

begin
end architecture;
